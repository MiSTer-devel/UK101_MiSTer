-- Copyright of the original ROM contents respectfully acknowleged

-- This file was created and maintaned by Grant Searle 2014
-- You are free to use this file in your own projects but must never charge for it nor use it without
-- acknowledgement.
-- Please ask permission from Grant Searle before republishing elsewhere.
-- If you use this file or any part of it, please add an acknowledgement to myself and
-- a link back to my main web site http://searle.hostei.com/grant/    
-- and to the UK101 page at http://searle.hostei.com/grant/uk101FPGA/index.html
--
-- Please check on the above web pages to see if there are any updates before using this file.
-- If for some reason the page is no longer available, please search for "Grant Searle"
-- on the internet to see if I have moved to another web hosting service.
--
-- Grant Searle
-- eMail address available on my main web page link above.

-- OSI character generator version - L.A. June 2017

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	use ieee.std_logic_unsigned.all;

ENTITY CharRomOSI IS

	PORT
	(
		address : in std_logic_vector(10 downto 0);
		q : out std_logic_vector(7 downto 0)
	);
END CharRomOSI;

architecture behavior of CharRomOSI is
type romtable is array (0 to 2047) of std_logic_vector(7 downto 0);
constant romdata : romtable :=
(
x"5A",x"7E",x"5A",x"18",x"18",x"5A",x"7E",x"5A",x"42",x"7E",x"5A",x"18",x"18",x"5A",x"7E",x"42",
x"81",x"42",x"24",x"24",x"24",x"24",x"42",x"81",x"81",x"42",x"3C",x"00",x"00",x"3C",x"42",x"81",
x"00",x"00",x"00",x"24",x"99",x"5A",x"FF",x"00",x"80",x"00",x"00",x"C0",x"C0",x"FC",x"FE",x"FC",
x"01",x"01",x"01",x"03",x"C7",x"FF",x"FF",x"7F",x"80",x"80",x"80",x"C0",x"E3",x"FF",x"FF",x"FE",
x"01",x"00",x"00",x"03",x"03",x"3F",x"7F",x"3F",x"00",x"00",x"FE",x"20",x"20",x"F8",x"E0",x"00",
x"00",x"00",x"18",x"FE",x"07",x"1F",x"1F",x"00",x"00",x"00",x"18",x"7F",x"E0",x"F8",x"F8",x"00",
x"00",x"00",x"7F",x"04",x"04",x"1F",x"07",x"00",x"18",x"3C",x"7E",x"FE",x"7E",x"3C",x"10",x"10",
x"00",x"00",x"18",x"3C",x"7E",x"7E",x"6A",x"7A",x"18",x"BC",x"FE",x"FF",x"B5",x"FF",x"B5",x"FD",
x"18",x"3C",x"5A",x"18",x"18",x"18",x"18",x"3C",x"F0",x"E0",x"F0",x"B8",x"1D",x"0E",x"04",x"08",
x"00",x"20",x"41",x"FF",x"FF",x"41",x"20",x"00",x"08",x"04",x"0E",x"1D",x"B8",x"F0",x"E0",x"F0",
x"3C",x"18",x"18",x"18",x"18",x"5A",x"3C",x"18",x"10",x"20",x"70",x"B8",x"1D",x"0F",x"07",x"0F",
x"00",x"04",x"82",x"FF",x"FF",x"82",x"04",x"00",x"0F",x"07",x"0F",x"1D",x"B8",x"70",x"20",x"10",
x"00",x"7C",x"52",x"7C",x"50",x"50",x"50",x"00",x"00",x"00",x"00",x"40",x"7E",x"02",x"00",x"00",
x"00",x"1C",x"14",x"14",x"3E",x"14",x"1C",x"00",x"00",x"1C",x"14",x"14",x"14",x"14",x"1C",x"00",
x"00",x"7E",x"40",x"48",x"4C",x"4E",x"0C",x"08",x"18",x"24",x"42",x"81",x"18",x"24",x"42",x"81",
x"00",x"7E",x"42",x"24",x"18",x"18",x"18",x"18",x"81",x"42",x"24",x"18",x"81",x"42",x"24",x"18",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"08",x"08",x"08",x"00",x"08",x"00",
x"14",x"14",x"14",x"00",x"00",x"00",x"00",x"00",x"14",x"14",x"3E",x"14",x"3E",x"14",x"14",x"00",
x"08",x"3C",x"0A",x"1C",x"28",x"1E",x"08",x"00",x"06",x"26",x"10",x"08",x"04",x"32",x"30",x"00",
x"04",x"0A",x"0A",x"04",x"2A",x"12",x"2C",x"00",x"08",x"08",x"08",x"00",x"00",x"00",x"00",x"00",
x"08",x"04",x"02",x"02",x"02",x"04",x"08",x"00",x"08",x"10",x"20",x"20",x"20",x"10",x"08",x"00",
x"08",x"2A",x"1C",x"08",x"1C",x"2A",x"08",x"00",x"00",x"08",x"08",x"3E",x"08",x"08",x"00",x"00",
x"00",x"00",x"00",x"00",x"08",x"08",x"04",x"00",x"00",x"00",x"00",x"3E",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"00",x"20",x"10",x"08",x"04",x"02",x"00",x"00",
x"1C",x"22",x"32",x"2A",x"26",x"22",x"1C",x"00",x"08",x"0C",x"08",x"08",x"08",x"08",x"1C",x"00",
x"1C",x"22",x"20",x"18",x"04",x"02",x"3E",x"00",x"3E",x"20",x"10",x"18",x"20",x"22",x"1C",x"00",
x"10",x"18",x"14",x"12",x"3E",x"10",x"10",x"00",x"3E",x"02",x"1E",x"20",x"20",x"22",x"1C",x"00",
x"38",x"04",x"02",x"1E",x"22",x"22",x"1C",x"00",x"3E",x"20",x"10",x"08",x"04",x"04",x"04",x"00",
x"1C",x"22",x"22",x"1C",x"22",x"22",x"1C",x"00",x"1C",x"22",x"22",x"3C",x"20",x"10",x"0E",x"00",
x"00",x"00",x"08",x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"08",x"00",x"08",x"08",x"04",x"00",
x"10",x"08",x"04",x"02",x"04",x"08",x"10",x"00",x"00",x"00",x"3E",x"00",x"3E",x"00",x"00",x"00",
x"04",x"08",x"10",x"20",x"10",x"08",x"04",x"00",x"1C",x"22",x"10",x"08",x"08",x"00",x"08",x"00",
x"1C",x"22",x"2A",x"3A",x"1A",x"02",x"3C",x"00",x"08",x"14",x"22",x"22",x"3E",x"22",x"22",x"00",
x"1E",x"22",x"22",x"1E",x"22",x"22",x"1E",x"00",x"1C",x"22",x"02",x"02",x"02",x"22",x"1C",x"00",
x"1E",x"22",x"22",x"22",x"22",x"22",x"1E",x"00",x"3E",x"02",x"02",x"1E",x"02",x"02",x"3E",x"00",
x"3E",x"02",x"02",x"1E",x"02",x"02",x"02",x"00",x"3C",x"02",x"02",x"02",x"32",x"22",x"3C",x"00",
x"22",x"22",x"22",x"3E",x"22",x"22",x"22",x"00",x"1C",x"08",x"08",x"08",x"08",x"08",x"1C",x"00",
x"20",x"20",x"20",x"20",x"20",x"22",x"1C",x"00",x"22",x"12",x"0A",x"06",x"0A",x"12",x"22",x"00",
x"02",x"02",x"02",x"02",x"02",x"02",x"3E",x"00",x"22",x"36",x"2A",x"2A",x"22",x"22",x"22",x"00",
x"22",x"22",x"26",x"2A",x"32",x"22",x"22",x"00",x"1C",x"22",x"22",x"22",x"22",x"22",x"1C",x"00",
x"1E",x"22",x"22",x"1E",x"02",x"02",x"02",x"00",x"1C",x"22",x"22",x"22",x"2A",x"12",x"2C",x"00",
x"1E",x"22",x"22",x"1E",x"0A",x"12",x"22",x"00",x"1C",x"22",x"02",x"1C",x"20",x"22",x"1C",x"00",
x"3E",x"08",x"08",x"08",x"08",x"08",x"08",x"00",x"22",x"22",x"22",x"22",x"22",x"22",x"1C",x"00",
x"22",x"22",x"22",x"22",x"22",x"14",x"08",x"00",x"22",x"22",x"22",x"2A",x"2A",x"36",x"22",x"00",
x"22",x"22",x"14",x"08",x"14",x"22",x"22",x"00",x"22",x"22",x"14",x"08",x"08",x"08",x"08",x"00",
x"3E",x"20",x"10",x"08",x"04",x"02",x"3E",x"00",x"3E",x"06",x"06",x"06",x"06",x"06",x"3E",x"00",
x"00",x"02",x"04",x"08",x"10",x"20",x"00",x"00",x"3E",x"30",x"30",x"30",x"30",x"30",x"3E",x"00",
x"00",x"00",x"08",x"14",x"22",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"3E",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2C",x"32",x"22",x"32",x"2C",x"00",
x"02",x"02",x"1A",x"26",x"22",x"26",x"1A",x"00",x"00",x"00",x"3C",x"02",x"02",x"02",x"3C",x"00",
x"20",x"20",x"2C",x"32",x"22",x"32",x"2C",x"00",x"00",x"00",x"1C",x"22",x"3E",x"02",x"1C",x"00",
x"10",x"08",x"08",x"1C",x"08",x"08",x"08",x"00",x"00",x"2C",x"32",x"22",x"32",x"2C",x"20",x"1C",
x"02",x"02",x"1E",x"22",x"22",x"22",x"22",x"00",x"00",x"08",x"00",x"0C",x"08",x"08",x"1C",x"00",
x"00",x"10",x"00",x"10",x"10",x"10",x"10",x"0C",x"02",x"22",x"12",x"0A",x"0E",x"12",x"22",x"00",
x"0C",x"08",x"08",x"08",x"08",x"08",x"1C",x"00",x"00",x"00",x"16",x"2A",x"2A",x"2A",x"2A",x"00",
x"00",x"00",x"1E",x"22",x"22",x"22",x"22",x"00",x"00",x"00",x"1C",x"22",x"22",x"22",x"1C",x"00",
x"00",x"1A",x"26",x"22",x"26",x"1A",x"02",x"02",x"00",x"2C",x"32",x"22",x"32",x"2C",x"20",x"20",
x"00",x"00",x"1A",x"06",x"02",x"02",x"02",x"00",x"00",x"00",x"3C",x"02",x"1C",x"20",x"1E",x"00",
x"00",x"08",x"3E",x"08",x"08",x"08",x"08",x"00",x"00",x"00",x"22",x"22",x"22",x"22",x"3C",x"00",
x"00",x"00",x"22",x"22",x"14",x"14",x"08",x"00",x"00",x"00",x"22",x"22",x"22",x"2A",x"14",x"00",
x"00",x"00",x"22",x"14",x"08",x"14",x"22",x"00",x"00",x"00",x"24",x"24",x"24",x"3C",x"20",x"1C",
x"00",x"00",x"3E",x"10",x"08",x"04",x"3E",x"00",x"30",x"08",x"08",x"04",x"08",x"08",x"30",x"00",
x"06",x"08",x"08",x"10",x"08",x"08",x"06",x"00",x"08",x"08",x"08",x"00",x"08",x"08",x"08",x"00",
x"00",x"08",x"00",x"3E",x"00",x"08",x"00",x"00",x"00",x"00",x"20",x"1C",x"02",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",
x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",
x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",
x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",
x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",
x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",
x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"F0",x"F0",x"F0",x"F0",
x"F0",x"F0",x"F0",x"F0",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",x"3C",x"3C",x"3C",x"3C",
x"3C",x"3C",x"3C",x"3C",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"00",x"00",
x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"FF",x"7F",x"3F",x"1F",x"0F",x"07",x"03",x"01",
x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",x"FF",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",
x"01",x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"FF",x"00",x"00",x"80",x"C2",x"EC",x"FF",x"FF",x"FF",
x"02",x"02",x"07",x"47",x"37",x"FF",x"7F",x"3F",x"40",x"40",x"E0",x"E2",x"EC",x"FF",x"FE",x"FC",
x"00",x"00",x"01",x"43",x"37",x"FF",x"FF",x"FF",x"55",x"AA",x"55",x"AA",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"55",x"AA",x"55",x"AA",x"05",x"0A",x"05",x"0A",x"05",x"0A",x"05",x"0A",
x"50",x"A0",x"50",x"A0",x"50",x"A0",x"50",x"A0",x"55",x"AA",x"55",x"AA",x"55",x"AA",x"55",x"AA",
x"81",x"42",x"24",x"18",x"18",x"24",x"42",x"81",x"80",x"40",x"20",x"10",x"08",x"04",x"02",x"01",
x"01",x"02",x"04",x"08",x"10",x"20",x"40",x"80",x"81",x"42",x"24",x"18",x"00",x"00",x"00",x"00",
x"80",x"40",x"20",x"10",x"10",x"20",x"40",x"80",x"00",x"00",x"00",x"00",x"18",x"24",x"42",x"81",
x"01",x"02",x"04",x"08",x"08",x"04",x"02",x"01",x"C0",x"30",x"0C",x"03",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"C0",x"30",x"0C",x"03",x"03",x"0C",x"30",x"C0",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"03",x"0C",x"30",x"C0",x"10",x"10",x"20",x"20",x"40",x"40",x"80",x"80",
x"01",x"01",x"02",x"02",x"04",x"04",x"08",x"08",x"80",x"80",x"40",x"40",x"20",x"20",x"10",x"10",
x"08",x"08",x"04",x"04",x"02",x"02",x"01",x"01",x"10",x"10",x"10",x"F0",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"F0",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"0F",x"08",x"08",x"08",
x"08",x"08",x"08",x"0F",x"00",x"00",x"00",x"00",x"FF",x"80",x"80",x"80",x"80",x"80",x"80",x"80",
x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"FF",
x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"07",x"8F",x"FF",x"F9",x"FF",x"00",x"00",
x"00",x"87",x"8F",x"FF",x"F0",x"FF",x"80",x"80",x"00",x"E1",x"F1",x"FF",x"0F",x"FF",x"01",x"01",
x"40",x"E0",x"F1",x"FF",x"9F",x"FF",x"00",x"00",x"18",x"18",x"18",x"FF",x"FF",x"00",x"00",x"00",
x"18",x"18",x"18",x"F8",x"F8",x"18",x"18",x"18",x"00",x"00",x"00",x"FF",x"FF",x"18",x"18",x"18",
x"18",x"18",x"18",x"1F",x"1F",x"18",x"18",x"18",x"18",x"18",x"18",x"FF",x"FF",x"18",x"18",x"18",
x"10",x"10",x"20",x"C0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"C0",x"20",x"10",x"10",
x"00",x"00",x"00",x"00",x"03",x"04",x"08",x"08",x"08",x"08",x"04",x"03",x"00",x"00",x"00",x"00",
x"C0",x"20",x"10",x"10",x"10",x"10",x"20",x"C0",x"03",x"04",x"08",x"08",x"08",x"08",x"04",x"03",
x"3C",x"42",x"81",x"81",x"81",x"81",x"42",x"3C",x"F0",x"0C",x"03",x"03",x"03",x"03",x"0C",x"F0",
x"0F",x"30",x"C0",x"C0",x"C0",x"C0",x"30",x"0F",x"66",x"FF",x"FF",x"FF",x"7E",x"3C",x"18",x"18",
x"3C",x"3C",x"18",x"42",x"E7",x"E7",x"18",x"3C",x"18",x"3C",x"7E",x"FF",x"FF",x"5A",x"18",x"3C",
x"18",x"3C",x"7E",x"FF",x"FF",x"7E",x"3C",x"18",x"E7",x"C3",x"81",x"00",x"00",x"81",x"C3",x"E7",
x"C0",x"F0",x"FC",x"FF",x"FF",x"FC",x"F0",x"C0",x"03",x"0F",x"3F",x"FF",x"FF",x"3F",x"0F",x"03",
x"18",x"18",x"3C",x"7E",x"FF",x"DB",x"18",x"3C",x"0C",x"1C",x"39",x"FF",x"FF",x"39",x"1C",x"0C",
x"3C",x"18",x"DB",x"FF",x"7E",x"3C",x"18",x"18",x"30",x"38",x"9C",x"FF",x"FF",x"9C",x"38",x"30",
x"00",x"00",x"00",x"08",x"1C",x"2A",x"08",x"14",x"00",x"00",x"40",x"48",x"3C",x"2A",x"18",x"14",
x"10",x"10",x"10",x"90",x"F0",x"F0",x"F8",x"F8",x"00",x"02",x"04",x"C8",x"F0",x"F0",x"F8",x"F8",
x"00",x"00",x"00",x"C0",x"FF",x"F0",x"F8",x"F8",x"08",x"08",x"08",x"09",x"0F",x"0F",x"1F",x"1F",
x"00",x"40",x"20",x"13",x"0F",x"0F",x"1F",x"1F",x"00",x"00",x"00",x"03",x"FF",x"0F",x"1F",x"1F",
x"00",x"10",x"10",x"54",x"7C",x"7C",x"7C",x"44",x"00",x"80",x"50",x"38",x"7C",x"3E",x"18",x"08",
x"00",x"1F",x"0E",x"7E",x"0E",x"1F",x"00",x"00",x"08",x"18",x"3E",x"7C",x"38",x"50",x"80",x"00",
x"44",x"7C",x"7C",x"7C",x"54",x"10",x"10",x"00",x"20",x"30",x"F8",x"7C",x"38",x"14",x"02",x"00",
x"00",x"F8",x"70",x"7E",x"70",x"F8",x"00",x"00",x"00",x"01",x"0A",x"1C",x"3E",x"7C",x"18",x"10"
);
begin
process (address)
begin
q <= romdata (to_integer(unsigned(address)));
end process;
end behavior;

