-- Copyright of the original ROM contents respectfully acknowleged

-- This file was created and maintaned by Grant Searle 2014
-- You are free to use this file in your own projects but must never charge for it nor use it without
-- acknowledgement.
-- Please ask permission from Grant Searle before republishing elsewhere.
-- If you use this file or any part of it, please add an acknowledgement to myself and
-- a link back to my main web site http://searle.hostei.com/grant/    
-- and to the UK101 page at http://searle.hostei.com/grant/uk101FPGA/index.html
--
-- Please check on the above web pages to see if there are any updates before using this file.
-- If for some reason the page is no longer available, please search for "Grant Searle"
-- on the internet to see if I have moved to another web hosting service.
--
-- Grant Searle
-- eMail address available on my main web page link above.

-- CEGMON C2/C4 version by Leslie Ayling
-- $FC00 block relocated to $F400
-- Register buf-fix included ($E1 -> $E4)

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	use ieee.std_logic_unsigned.all;

ENTITY WemonRom IS

	PORT
	(
		address : in std_logic_vector(11 downto 0);
		q : out std_logic_vector(7 downto 0)
	);
END WemonRom;

architecture behavior of WemonRom is
type romtable is array (0 to 4095) of std_logic_vector(7 downto 0);
constant romdata : romtable :=
(
x"A2",x"28",x"9A",x"D8",x"A9",x"7F",x"8D",x"2D",
x"02",x"A9",x"06",x"8D",x"40",x"02",x"A9",x"00",
x"8D",x"03",x"02",x"8D",x"4F",x"02",x"8D",x"05",
x"02",x"8D",x"22",x"02",x"8D",x"27",x"02",x"8D",
x"23",x"02",x"8D",x"24",x"02",x"8D",x"26",x"02",
x"8D",x"12",x"02",x"8D",x"04",x"02",x"8D",x"4E",
x"02",x"8D",x"4B",x"02",x"8D",x"06",x"02",x"A9",
x"98",x"8D",x"4C",x"02",x"20",x"EF",x"FE",x"A0",
x"09",x"B9",x"78",x"F7",x"99",x"18",x"02",x"88",
x"10",x"F7",x"A9",x"00",x"85",x"F6",x"85",x"E0",
x"85",x"D6",x"20",x"94",x"F0",x"A9",x"A1",x"8D",
x"2C",x"02",x"20",x"A2",x"F0",x"A2",x"00",x"20",
x"82",x"F7",x"20",x"69",x"F3",x"29",x"5F",x"C9",
x"4D",x"D0",x"0A",x"A9",x"F0",x"48",x"A9",x"5E",
x"48",x"08",x"4C",x"55",x"F8",x"C9",x"43",x"D0",
x"03",x"4C",x"11",x"BD",x"C9",x"57",x"D0",x"03",
x"4C",x"74",x"A2",x"C9",x"44",x"D0",x"03",x"6C",
x"4B",x"02",x"C9",x"55",x"D0",x"D4",x"20",x"29",
x"02",x"4C",x"62",x"F0",x"A9",x"03",x"8D",x"00",
x"E0",x"A9",x"11",x"8D",x"00",x"E0",x"8D",x"4F",
x"02",x"60",x"A9",x"60",x"A0",x"00",x"8D",x"01",
x"02",x"99",x"00",x"D3",x"99",x"00",x"D2",x"99",
x"00",x"D1",x"99",x"00",x"D0",x"C8",x"D0",x"F1",
x"A9",x"D0",x"8D",x"25",x"02",x"85",x"F7",x"A0",
x"4B",x"8C",x"00",x"02",x"D0",x"48",x"A9",x"00",
x"85",x"F6",x"AD",x"25",x"02",x"85",x"F7",x"AC",
x"00",x"02",x"60",x"8D",x"02",x"02",x"48",x"8A",
x"48",x"98",x"48",x"20",x"C6",x"F0",x"20",x"ED",
x"F0",x"20",x"29",x"F2",x"4C",x"37",x"F2",x"AD",
x"01",x"02",x"91",x"F6",x"60",x"AD",x"02",x"02",
x"C9",x"0D",x"D0",x"30",x"20",x"5C",x"F2",x"C0",
x"CA",x"F0",x"09",x"20",x"88",x"F1",x"A9",x"60",
x"D1",x"F6",x"F0",x"07",x"20",x"75",x"F1",x"A9",
x"60",x"91",x"F6",x"C8",x"C6",x"D6",x"A9",x"00",
x"85",x"F6",x"8D",x"26",x"02",x"8D",x"27",x"02",
x"8D",x"22",x"02",x"8D",x"23",x"02",x"A9",x"A1",
x"8D",x"2C",x"02",x"60",x"C9",x"22",x"D0",x"03",
x"20",x"01",x"F5",x"C9",x"20",x"90",x"17",x"C9",
x"3F",x"D0",x"10",x"20",x"4A",x"F2",x"D0",x"09",
x"A9",x"FF",x"C5",x"88",x"F0",x"03",x"8D",x"04",
x"02",x"A9",x"3F",x"4C",x"EF",x"F1",x"C9",x"0E",
x"F0",x"0B",x"2C",x"26",x"02",x"10",x"06",x"20",
x"D6",x"F1",x"4C",x"EF",x"F1",x"C9",x"08",x"D0",
x"18",x"88",x"20",x"4A",x"F2",x"B0",x"11",x"20",
x"3F",x"F2",x"B0",x"09",x"A9",x"D0",x"85",x"F3",
x"A0",x"7B",x"4C",x"B0",x"F2",x"20",x"50",x"F2",
x"60",x"C9",x"0A",x"D0",x"21",x"A5",x"D6",x"D0",
x"18",x"C0",x"CA",x"90",x"0B",x"A9",x"D3",x"C5",
x"F7",x"D0",x"05",x"85",x"F3",x"4C",x"65",x"F2",
x"98",x"18",x"69",x"40",x"A8",x"90",x"02",x"E6",
x"F7",x"A9",x"00",x"85",x"D6",x"60",x"C9",x"09",
x"F0",x"57",x"C9",x"1A",x"D0",x"1B",x"C0",x"8B",
x"B0",x"0B",x"A9",x"D0",x"C5",x"F7",x"D0",x"05",
x"85",x"F3",x"4C",x"B0",x"F2",x"48",x"98",x"38",
x"E9",x"40",x"A8",x"B0",x"02",x"C6",x"F7",x"68",
x"60",x"C9",x"0C",x"D0",x"03",x"4C",x"A2",x"F0",
x"C9",x"01",x"D0",x"03",x"4C",x"B8",x"F0",x"C9",
x"0E",x"D0",x"03",x"4C",x"AB",x"F6",x"C9",x"1E",
x"D0",x"03",x"4C",x"E7",x"F5",x"60",x"85",x"EC",
x"98",x"48",x"20",x"CB",x"F5",x"20",x"D4",x"F5",
x"C9",x"FF",x"F0",x"06",x"20",x"C2",x"F5",x"20",
x"E2",x"F5",x"68",x"A8",x"A5",x"EC",x"60",x"91",
x"F6",x"C8",x"20",x"1A",x"F2",x"90",x"0D",x"20",
x"0C",x"F2",x"B0",x"09",x"20",x"22",x"F2",x"A9",
x"20",x"91",x"F6",x"C8",x"60",x"A0",x"CA",x"20",
x"65",x"F2",x"D0",x"F3",x"48",x"98",x"C9",x"FB",
x"B0",x"02",x"68",x"60",x"A5",x"F7",x"C9",x"D3",
x"68",x"60",x"48",x"98",x"29",x"3F",x"C9",x"3B",
x"68",x"60",x"20",x"5C",x"F2",x"20",x"88",x"F1",
x"60",x"B1",x"F6",x"8D",x"01",x"02",x"A5",x"F7",
x"8D",x"25",x"02",x"8C",x"00",x"02",x"60",x"68",
x"A8",x"68",x"AA",x"68",x"4C",x"6C",x"FF",x"C0",
x"4B",x"B0",x"06",x"48",x"A5",x"F7",x"C9",x"D1",
x"68",x"60",x"98",x"29",x"3F",x"C9",x"0B",x"60",
x"48",x"98",x"38",x"E9",x"10",x"A8",x"B0",x"02",
x"C6",x"F7",x"68",x"60",x"48",x"98",x"29",x"C0",
x"09",x"0A",x"A8",x"68",x"60",x"20",x"8A",x"F2",
x"AC",x"06",x"02",x"F0",x"03",x"20",x"0D",x"F7",
x"20",x"3E",x"F8",x"D0",x"12",x"A9",x"03",x"85",
x"E5",x"A0",x"C0",x"20",x"0D",x"F7",x"20",x"3E",
x"F8",x"D0",x"04",x"C6",x"E5",x"D0",x"F4",x"4C",
x"C6",x"F0",x"20",x"2E",x"F2",x"A0",x"40",x"A2",
x"CF",x"A9",x"40",x"85",x"F8",x"E8",x"86",x"F9",
x"86",x"F7",x"B1",x"F8",x"91",x"F6",x"C8",x"D0",
x"F9",x"E0",x"D3",x"D0",x"F0",x"A9",x"60",x"88",
x"91",x"F6",x"88",x"C0",x"C0",x"D0",x"F9",x"60",
x"20",x"B5",x"F2",x"30",x"D2",x"20",x"2E",x"F2",
x"98",x"29",x"C0",x"85",x"F4",x"A0",x"BF",x"A9",
x"40",x"85",x"F8",x"A2",x"D4",x"CA",x"86",x"F7",
x"86",x"F9",x"B1",x"F6",x"91",x"F8",x"C4",x"F4",
x"D0",x"04",x"E4",x"F3",x"F0",x"07",x"88",x"C0",
x"FF",x"D0",x"EF",x"F0",x"E8",x"A9",x"3F",x"85",
x"F8",x"AD",x"00",x"02",x"29",x"C0",x"A8",x"A9",
x"60",x"91",x"F8",x"C6",x"F8",x"10",x"FA",x"60",
x"AD",x"04",x"02",x"F0",x"16",x"30",x"08",x"A9",
x"00",x"8D",x"04",x"02",x"4C",x"74",x"A2",x"A9",
x"00",x"C5",x"8C",x"D0",x"03",x"4C",x"D2",x"F4",
x"8D",x"04",x"02",x"98",x"48",x"8A",x"48",x"20",
x"69",x"F3",x"C9",x"0D",x"F0",x"17",x"C9",x"0E",
x"F0",x"09",x"2C",x"26",x"02",x"30",x"1E",x"C9",
x"20",x"B0",x"1A",x"2C",x"27",x"02",x"30",x"27",
x"CE",x"27",x"02",x"D0",x"22",x"20",x"C6",x"F0",
x"AD",x"01",x"02",x"91",x"F6",x"2C",x"27",x"02",
x"10",x"1E",x"4C",x"7D",x"F5",x"68",x"48",x"AA",
x"AD",x"13",x"02",x"95",x"13",x"86",x"DF",x"E8",
x"68",x"8A",x"48",x"E0",x"47",x"F0",x"09",x"AD",
x"13",x"02",x"20",x"D3",x"F0",x"4C",x"0F",x"F3",
x"68",x"AA",x"68",x"A8",x"86",x"F8",x"BA",x"E8",
x"E8",x"E8",x"E8",x"9A",x"A6",x"F8",x"4C",x"66",
x"A8",x"98",x"48",x"8A",x"48",x"A9",x"02",x"20",
x"16",x"F7",x"20",x"1E",x"F7",x"D0",x"1A",x"0A",
x"D0",x"F5",x"A9",x"01",x"20",x"16",x"F7",x"20",
x"27",x"F7",x"85",x"EC",x"29",x"FE",x"C9",x"44",
x"D0",x"3A",x"A9",x"FF",x"8D",x"24",x"02",x"D0",
x"DC",x"4A",x"20",x"FE",x"F3",x"98",x"8D",x"13",
x"02",x"0A",x"0A",x"0A",x"38",x"ED",x"13",x"02",
x"8D",x"13",x"02",x"8A",x"4A",x"20",x"FE",x"F3",
x"D0",x"1A",x"98",x"18",x"6D",x"13",x"02",x"A8",
x"B9",x"8D",x"FE",x"CD",x"15",x"02",x"D0",x"3B",
x"CE",x"14",x"02",x"F0",x"48",x"A0",x"05",x"20",
x"0D",x"F7",x"F0",x"A9",x"24",x"D7",x"30",x"21",
x"C6",x"D7",x"D0",x"22",x"CE",x"40",x"02",x"D0",
x"18",x"20",x"C6",x"F0",x"AD",x"01",x"02",x"D1",
x"F6",x"F0",x"04",x"91",x"F6",x"D0",x"05",x"AD",
x"2C",x"02",x"91",x"F6",x"A9",x"06",x"8D",x"40",
x"02",x"AD",x"2D",x"02",x"85",x"D7",x"A9",x"00",
x"8D",x"16",x"02",x"8D",x"15",x"02",x"A9",x"02",
x"8D",x"14",x"02",x"4C",x"6D",x"F3",x"A0",x"08",
x"88",x"0A",x"90",x"FC",x"60",x"48",x"98",x"48",
x"20",x"C6",x"F0",x"AD",x"01",x"02",x"91",x"F6",
x"68",x"A8",x"68",x"2C",x"24",x"02",x"10",x"03",
x"4C",x"17",x"F5",x"A2",x"96",x"CD",x"16",x"02",
x"D0",x"02",x"A2",x"14",x"8E",x"14",x"02",x"8D",
x"16",x"02",x"A5",x"EC",x"29",x"40",x"D0",x"36",
x"A5",x"EC",x"4A",x"29",x"03",x"D0",x"12",x"90",
x"05",x"AD",x"15",x"02",x"D0",x"5E",x"AD",x"15",
x"02",x"C9",x"41",x"90",x"57",x"09",x"20",x"D0",
x"53",x"AD",x"15",x"02",x"C9",x"41",x"B0",x"4C",
x"C9",x"20",x"F0",x"48",x"C9",x"0D",x"F0",x"44",
x"C9",x"30",x"F0",x"40",x"B0",x"04",x"09",x"10",
x"D0",x"3A",x"29",x"2F",x"D0",x"36",x"AD",x"15",
x"02",x"29",x"1F",x"C9",x"10",x"D0",x"08",x"A9",
x"FF",x"4D",x"4E",x"02",x"4C",x"6D",x"F3",x"C9",
x"11",x"D0",x"05",x"20",x"01",x"F5",x"D0",x"10",
x"C9",x"14",x"D0",x"05",x"20",x"2D",x"F7",x"D0",
x"07",x"C9",x"04",x"D0",x"06",x"20",x"50",x"F5",
x"4C",x"6D",x"F3",x"C9",x"05",x"D0",x"05",x"20",
x"A7",x"F4",x"30",x"F4",x"8D",x"13",x"02",x"68",
x"AA",x"68",x"A8",x"AD",x"13",x"02",x"60",x"A2",
x"03",x"BD",x"B2",x"F4",x"95",x"C5",x"CA",x"10",
x"F8",x"60",x"4C",x"B6",x"F4",x"EA",x"08",x"48",
x"A5",x"C4",x"D0",x"11",x"A6",x"DF",x"D0",x"0D",
x"68",x"48",x"C9",x"41",x"90",x"07",x"C9",x"5B",
x"B0",x"03",x"20",x"48",x"02",x"68",x"28",x"4C",
x"F7",x"BC",x"A5",x"88",x"A4",x"87",x"20",x"C1",
x"AF",x"20",x"6E",x"B9",x"A2",x"00",x"A0",x"39",
x"B9",x"8E",x"F7",x"F0",x"06",x"95",x"13",x"C8",
x"E8",x"D0",x"F5",x"A0",x"00",x"B9",x"01",x"01",
x"F0",x"07",x"9D",x"13",x"00",x"C8",x"E8",x"D0",
x"F4",x"A9",x"7F",x"8D",x"04",x"02",x"4C",x"5C",
x"F3",x"48",x"A9",x"FF",x"4D",x"26",x"02",x"8D",
x"26",x"02",x"10",x"04",x"A9",x"17",x"D0",x"02",
x"A9",x"A1",x"8D",x"2C",x"02",x"68",x"60",x"B9",
x"BE",x"FE",x"A8",x"BA",x"BD",x"05",x"01",x"AA",
x"B9",x"84",x"A0",x"48",x"29",x"7F",x"20",x"69",
x"FF",x"68",x"30",x"06",x"95",x"13",x"C8",x"E8",
x"D0",x"EE",x"29",x"7F",x"95",x"13",x"E8",x"C9",
x"24",x"D0",x"08",x"A9",x"28",x"20",x"69",x"FF",
x"95",x"13",x"E8",x"8A",x"BA",x"9D",x"05",x"01",
x"A9",x"00",x"8D",x"24",x"02",x"4C",x"6D",x"F3",
x"20",x"C6",x"F0",x"AD",x"25",x"02",x"C0",x"CB",
x"90",x"05",x"C9",x"D3",x"90",x"01",x"60",x"85",
x"F3",x"20",x"B8",x"F2",x"A9",x"60",x"8D",x"01",
x"02",x"D0",x"F3",x"20",x"5C",x"F2",x"B1",x"F6",
x"C9",x"60",x"F0",x"08",x"20",x"3F",x"F2",x"90",
x"03",x"20",x"AD",x"F1",x"60",x"A2",x"00",x"20",
x"6B",x"F5",x"C8",x"20",x"1A",x"F2",x"90",x"0D",
x"E0",x"31",x"B0",x"2E",x"20",x"0C",x"F2",x"B0",
x"29",x"20",x"22",x"F2",x"C8",x"B1",x"F6",x"C9",
x"60",x"F0",x"1F",x"85",x"EC",x"98",x"48",x"20",
x"C2",x"F5",x"20",x"D4",x"F5",x"C9",x"FF",x"F0",
x"06",x"20",x"CB",x"F5",x"20",x"E2",x"F5",x"68",
x"A8",x"A5",x"EC",x"95",x"13",x"E8",x"E0",x"47",
x"D0",x"C8",x"8A",x"BA",x"9D",x"01",x"01",x"4C",
x"58",x"F3",x"A9",x"D7",x"85",x"FE",x"A9",x"FF",
x"85",x"FF",x"60",x"A9",x"49",x"85",x"FE",x"A9",
x"FF",x"85",x"FF",x"60",x"A5",x"EC",x"A0",x"06",
x"D1",x"FE",x"F0",x"05",x"88",x"10",x"F9",x"A9",
x"FF",x"60",x"B1",x"FE",x"85",x"EC",x"60",x"2C",
x"23",x"02",x"30",x"41",x"20",x"6B",x"F5",x"A2",
x"00",x"C8",x"A9",x"60",x"D1",x"F6",x"D0",x"0D",
x"E0",x"00",x"F0",x"31",x"E0",x"47",x"90",x"32",
x"CE",x"23",x"02",x"D0",x"28",x"E0",x"47",x"B0",
x"F7",x"E8",x"C8",x"20",x"1A",x"F2",x"90",x"E2",
x"E0",x"31",x"B0",x"19",x"20",x"0C",x"F2",x"B0",
x"18",x"20",x"22",x"F2",x"B1",x"F6",x"C8",x"C9",
x"60",x"F0",x"05",x"CE",x"22",x"02",x"D0",x"CA",
x"20",x"50",x"F2",x"D0",x"05",x"20",x"C6",x"F0",
x"60",x"88",x"A5",x"F7",x"48",x"98",x"48",x"B1",
x"F6",x"48",x"C8",x"20",x"1A",x"F2",x"90",x"44",
x"2C",x"22",x"02",x"30",x"20",x"CE",x"22",x"02",
x"20",x"0C",x"F2",x"B0",x"1E",x"20",x"22",x"F2",
x"A5",x"F7",x"85",x"F3",x"48",x"98",x"48",x"20",
x"B8",x"F2",x"68",x"A8",x"68",x"85",x"F7",x"A9",
x"20",x"91",x"F6",x"D0",x"03",x"20",x"22",x"F2",
x"C8",x"D0",x"19",x"AD",x"00",x"02",x"38",x"E9",
x"40",x"8D",x"00",x"02",x"BA",x"A9",x"BA",x"9D",
x"02",x"01",x"20",x"8D",x"F2",x"A0",x"CA",x"A9",
x"20",x"91",x"F6",x"C8",x"68",x"91",x"F6",x"68",
x"A8",x"68",x"85",x"F7",x"CC",x"00",x"02",x"F0",
x"0B",x"88",x"20",x"4A",x"F2",x"B0",x"9B",x"20",
x"50",x"F2",x"D0",x"96",x"AD",x"01",x"02",x"C8",
x"91",x"F6",x"A9",x"20",x"88",x"91",x"F6",x"8D",
x"01",x"02",x"60",x"20",x"E7",x"F0",x"20",x"6B",
x"F5",x"C8",x"CC",x"00",x"02",x"F0",x"3F",x"20",
x"C6",x"F0",x"CE",x"00",x"02",x"AD",x"00",x"02",
x"29",x"3F",x"C9",x"0A",x"D0",x"0E",x"AD",x"00",
x"02",x"38",x"E9",x"10",x"8D",x"00",x"02",x"B0",
x"03",x"CE",x"25",x"02",x"A5",x"F7",x"48",x"98",
x"48",x"B1",x"F6",x"48",x"88",x"20",x"4A",x"F2",
x"B0",x"08",x"20",x"3F",x"F2",x"90",x"21",x"20",
x"50",x"F2",x"68",x"91",x"F6",x"C9",x"60",x"D0",
x"06",x"68",x"68",x"20",x"C6",x"F0",x"60",x"68",
x"A8",x"68",x"85",x"F7",x"C8",x"20",x"1A",x"F2",
x"90",x"D2",x"20",x"22",x"F2",x"C8",x"D0",x"CC",
x"68",x"68",x"4C",x"2B",x"F2",x"A2",x"C8",x"CA",
x"D0",x"FD",x"88",x"D0",x"F8",x"60",x"49",x"FF",
x"8D",x"00",x"DF",x"49",x"FF",x"60",x"48",x"20",
x"27",x"F7",x"AA",x"68",x"CA",x"E8",x"60",x"AD",
x"00",x"DF",x"49",x"FF",x"60",x"2C",x"4F",x"02",
x"30",x"0B",x"A9",x"51",x"8D",x"00",x"E0",x"0A",
x"8D",x"4F",x"02",x"D0",x"08",x"A9",x"11",x"8D",
x"00",x"E0",x"8D",x"4F",x"02",x"60",x"A9",x"00",
x"8D",x"05",x"02",x"8D",x"03",x"02",x"85",x"E0",
x"20",x"3D",x"F7",x"60",x"A2",x"06",x"A9",x"00",
x"20",x"5F",x"F7",x"CA",x"D0",x"FA",x"60",x"48",
x"20",x"3E",x"F8",x"F0",x"0E",x"68",x"48",x"AD",
x"00",x"E0",x"4A",x"4A",x"90",x"F9",x"68",x"8D",
x"01",x"E0",x"60",x"20",x"46",x"F7",x"68",x"60",
x"BA",x"FF",x"D3",x"F0",x"9A",x"FF",x"8B",x"FF",
x"96",x"FF",x"BD",x"8E",x"F7",x"F0",x"06",x"20",
x"69",x"FF",x"E8",x"D0",x"F5",x"60",x"57",x"45",
x"4D",x"4F",x"4E",x"20",x"28",x"43",x"29",x"31",
x"39",x"38",x"31",x"2E",x"0D",x"0A",x"4D",x"2F",
x"43",x"2F",x"57",x"2F",x"44",x"2F",x"55",x"20",
x"3F",x"00",x"0D",x"0A",x"46",x"4F",x"55",x"4E",
x"44",x"20",x"00",x"0D",x"0A",x"4C",x"4F",x"41",
x"44",x"49",x"4E",x"47",x"00",x"0D",x"0A",x"53",
x"41",x"56",x"49",x"4E",x"47",x"20",x"00",x"4C",
x"49",x"53",x"54",x"00",x"C9",x"30",x"30",x"12",
x"C9",x"3A",x"30",x"0B",x"C9",x"41",x"30",x"0A",
x"C9",x"47",x"10",x"06",x"38",x"E9",x"07",x"29",
x"0F",x"60",x"A9",x"80",x"60",x"A2",x"03",x"20",
x"F6",x"F7",x"E0",x"02",x"D0",x"04",x"20",x"13",
x"F8",x"CA",x"CA",x"10",x"F2",x"60",x"B5",x"FA",
x"4A",x"4A",x"4A",x"4A",x"20",x"18",x"F8",x"B5",
x"FA",x"4C",x"18",x"F8",x"A9",x"0D",x"20",x"69",
x"FF",x"A9",x"0A",x"4C",x"69",x"FF",x"A9",x"20",
x"20",x"69",x"FF",x"A9",x"20",x"4C",x"69",x"FF",
x"29",x"0F",x"09",x"30",x"C9",x"3A",x"30",x"03",
x"18",x"69",x"07",x"D0",x"F0",x"A0",x"04",x"0A",
x"0A",x"0A",x"0A",x"2A",x"36",x"FA",x"36",x"FB",
x"88",x"D0",x"F8",x"60",x"A5",x"E0",x"F0",x"03",
x"4C",x"C2",x"FF",x"4C",x"69",x"F3",x"A9",x"FD",
x"8D",x"00",x"DF",x"A9",x"10",x"2C",x"00",x"DF",
x"60",x"8D",x"45",x"02",x"68",x"48",x"29",x"10",
x"D0",x"06",x"6C",x"32",x"02",x"8D",x"45",x"02",
x"8E",x"46",x"02",x"8C",x"47",x"02",x"68",x"8D",
x"43",x"02",x"68",x"38",x"E9",x"01",x"8D",x"42",
x"02",x"68",x"E9",x"00",x"8D",x"41",x"02",x"BA",
x"8E",x"44",x"02",x"A2",x"28",x"9A",x"D8",x"20",
x"A2",x"F0",x"20",x"69",x"F9",x"20",x"B8",x"F0",
x"20",x"DD",x"F2",x"20",x"69",x"F3",x"85",x"EF",
x"20",x"69",x"FF",x"20",x"13",x"F8",x"A5",x"EF",
x"C9",x"52",x"D0",x"09",x"20",x"B8",x"F0",x"20",
x"F5",x"F8",x"4C",x"01",x"F9",x"C9",x"53",x"D0",
x"03",x"4C",x"BF",x"FC",x"C9",x"4C",x"D0",x"03",
x"4C",x"FD",x"FC",x"20",x"D5",x"F9",x"A5",x"EF",
x"C9",x"4D",x"D0",x"17",x"A5",x"E1",x"F0",x"0D",
x"C9",x"03",x"F0",x"06",x"20",x"F0",x"F8",x"4C",
x"AB",x"F8",x"4C",x"5F",x"FA",x"20",x"04",x"F8",
x"4C",x"07",x"FE",x"C9",x"46",x"D0",x"03",x"4C",
x"A0",x"FA",x"C9",x"42",x"D0",x"03",x"4C",x"EC",
x"FA",x"C9",x"56",x"D0",x"03",x"4C",x"21",x"FA",
x"C9",x"47",x"D0",x"03",x"4C",x"BA",x"FA",x"20",
x"29",x"02",x"20",x"04",x"F8",x"4C",x"83",x"F8",
x"A9",x"0D",x"20",x"69",x"FF",x"20",x"DD",x"F2",
x"A5",x"EF",x"20",x"69",x"FF",x"20",x"13",x"F8",
x"60",x"A9",x"00",x"85",x"EA",x"20",x"1B",x"FA",
x"D0",x"06",x"20",x"69",x"FF",x"4C",x"7A",x"F8",
x"C9",x"30",x"B0",x"12",x"C9",x"20",x"F0",x"08",
x"C9",x"08",x"F0",x"04",x"C9",x"18",x"D0",x"03",
x"20",x"69",x"FF",x"4C",x"01",x"F9",x"85",x"E9",
x"A5",x"EA",x"D0",x"14",x"AD",x"00",x"02",x"38",
x"E9",x"40",x"A0",x"06",x"D9",x"CD",x"F9",x"F0",
x"05",x"88",x"10",x"F8",x"30",x"C3",x"84",x"EB",
x"A5",x"E9",x"20",x"CC",x"F7",x"30",x"BE",x"48",
x"A5",x"E9",x"20",x"69",x"FF",x"68",x"A6",x"EA",
x"D0",x"04",x"A2",x"02",x"86",x"EA",x"A2",x"00",
x"20",x"25",x"F8",x"C6",x"EA",x"D0",x"A6",x"A6",
x"EB",x"A5",x"FA",x"9D",x"41",x"02",x"4C",x"01",
x"F9",x"A0",x"0C",x"A2",x"00",x"BD",x"A8",x"F9",
x"F0",x"07",x"99",x"00",x"D0",x"C8",x"E8",x"D0",
x"F4",x"A2",x"00",x"BC",x"CD",x"F9",x"F0",x"06",
x"20",x"87",x"F9",x"E8",x"D0",x"F5",x"60",x"BD",
x"41",x"02",x"4A",x"4A",x"4A",x"4A",x"20",x"99",
x"F9",x"BD",x"41",x"02",x"C8",x"20",x"99",x"F9",
x"60",x"29",x"0F",x"09",x"30",x"C9",x"3A",x"30",
x"03",x"18",x"69",x"07",x"99",x"00",x"D0",x"60",
x"50",x"43",x"20",x"20",x"20",x"20",x"20",x"20",
x"46",x"52",x"20",x"20",x"20",x"20",x"53",x"50",
x"20",x"20",x"20",x"20",x"41",x"43",x"43",x"20",
x"20",x"20",x"20",x"58",x"52",x"20",x"20",x"20",
x"20",x"59",x"52",x"20",x"00",x"0F",x"11",x"17",
x"1D",x"24",x"2A",x"30",x"00",x"A2",x"05",x"A9",
x"00",x"95",x"FA",x"CA",x"10",x"FB",x"E8",x"86",
x"E1",x"86",x"E3",x"20",x"1B",x"FA",x"F0",x"32",
x"E6",x"E1",x"D0",x"05",x"20",x"1B",x"FA",x"F0",
x"29",x"C9",x"2D",x"F0",x"15",x"85",x"E4",x"20",
x"CC",x"F7",x"30",x"F0",x"48",x"A5",x"E4",x"20",
x"69",x"FF",x"68",x"A6",x"E3",x"20",x"25",x"F8",
x"F0",x"E2",x"20",x"69",x"FF",x"A5",x"E1",x"0A",
x"85",x"E3",x"E6",x"E1",x"A6",x"E1",x"E0",x"04",
x"D0",x"D2",x"60",x"20",x"69",x"F3",x"C9",x"0D",
x"60",x"20",x"38",x"FD",x"A6",x"E1",x"E0",x"02",
x"F0",x"06",x"20",x"F0",x"F8",x"4C",x"21",x"FA",
x"A2",x"07",x"86",x"E4",x"20",x"04",x"F8",x"A2",
x"03",x"20",x"F6",x"F7",x"CA",x"20",x"F6",x"F7",
x"20",x"13",x"F8",x"A0",x"00",x"B1",x"FC",x"85",
x"FA",x"A2",x"00",x"20",x"F6",x"F7",x"20",x"13",
x"F8",x"20",x"33",x"FF",x"B0",x"06",x"C6",x"E4",
x"10",x"E9",x"30",x"D4",x"4C",x"EA",x"F8",x"20",
x"04",x"F8",x"A2",x"00",x"86",x"DE",x"86",x"DF",
x"A0",x"00",x"A5",x"FA",x"D1",x"FC",x"D0",x"17",
x"20",x"E5",x"F7",x"20",x"04",x"F8",x"F8",x"18",
x"AD",x"DE",x"00",x"69",x"01",x"85",x"DE",x"90",
x"06",x"A5",x"DF",x"69",x"00",x"85",x"DF",x"D8",
x"20",x"33",x"FF",x"90",x"DB",x"A5",x"DE",x"85",
x"FA",x"A5",x"DF",x"85",x"FB",x"A2",x"01",x"20",
x"F6",x"F7",x"CA",x"10",x"FA",x"4C",x"EA",x"F8",
x"A5",x"E1",x"C9",x"03",x"F0",x"06",x"20",x"F0",
x"F8",x"4C",x"A0",x"FA",x"A0",x"00",x"A5",x"FA",
x"91",x"FC",x"20",x"33",x"FF",x"90",x"F5",x"4C",
x"EA",x"F8",x"A5",x"E1",x"F0",x"0A",x"A5",x"FA",
x"8D",x"42",x"02",x"A5",x"FB",x"8D",x"41",x"02",
x"AD",x"41",x"02",x"48",x"AD",x"42",x"02",x"8D",
x"41",x"02",x"68",x"8D",x"42",x"02",x"AE",x"44",
x"02",x"9A",x"AE",x"46",x"02",x"AC",x"47",x"02",
x"AD",x"43",x"02",x"48",x"AD",x"45",x"02",x"28",
x"58",x"6C",x"41",x"02",x"A5",x"E1",x"C9",x"03",
x"F0",x"06",x"20",x"F0",x"F8",x"4C",x"EC",x"FA",
x"A5",x"FD",x"C5",x"FB",x"90",x"1A",x"A5",x"FC",
x"C5",x"FA",x"90",x"14",x"A0",x"00",x"B1",x"FC",
x"91",x"FA",x"E6",x"FA",x"D0",x"02",x"E6",x"FB",
x"20",x"33",x"FF",x"90",x"F1",x"4C",x"EA",x"F8",
x"20",x"42",x"FD",x"A2",x"00",x"20",x"42",x"FB",
x"A2",x"01",x"B5",x"F8",x"49",x"FF",x"95",x"F8",
x"CA",x"10",x"F7",x"C6",x"FF",x"C6",x"FB",x"A0",
x"FF",x"B1",x"FE",x"91",x"FA",x"E6",x"F8",x"D0",
x"04",x"E6",x"F9",x"F0",x"D8",x"88",x"D0",x"F1",
x"F0",x"E9",x"A5",x"F8",x"18",x"65",x"FA",x"95",
x"FA",x"A5",x"F9",x"65",x"FB",x"95",x"FB",x"60",
x"48",x"98",x"48",x"8A",x"48",x"20",x"96",x"FC",
x"20",x"B2",x"FC",x"20",x"CB",x"FB",x"B1",x"FC",
x"D0",x"0F",x"CA",x"D0",x"0E",x"20",x"5F",x"F7",
x"20",x"46",x"F7",x"68",x"AA",x"68",x"A8",x"68",
x"60",x"A2",x"03",x"20",x"5F",x"F7",x"20",x"C4",
x"FB",x"D0",x"E3",x"A9",x"14",x"85",x"DD",x"A0",
x"FF",x"20",x"0D",x"F7",x"C6",x"DD",x"D0",x"F7",
x"60",x"20",x"96",x"FC",x"20",x"D6",x"FB",x"A6",
x"E2",x"D0",x"04",x"CE",x"03",x"02",x"60",x"20",
x"CB",x"FB",x"20",x"C7",x"FF",x"D0",x"1C",x"CA",
x"D0",x"1B",x"91",x"FC",x"20",x"C4",x"FB",x"A5",
x"FC",x"85",x"7B",x"A5",x"FD",x"85",x"7C",x"A9",
x"01",x"85",x"79",x"A9",x"03",x"85",x"7A",x"20",
x"46",x"F7",x"60",x"A2",x"03",x"91",x"FC",x"20",
x"C4",x"FB",x"D0",x"D6",x"E6",x"FC",x"D0",x"02",
x"E6",x"FD",x"60",x"A9",x"03",x"85",x"FD",x"AA",
x"A9",x"00",x"85",x"FC",x"A8",x"60",x"20",x"32",
x"F7",x"A6",x"E0",x"D0",x"04",x"A6",x"E2",x"F0",
x"17",x"20",x"13",x"FC",x"20",x"3F",x"FC",x"A2",
x"1C",x"20",x"82",x"F7",x"20",x"23",x"FF",x"A6",
x"E2",x"F0",x"05",x"20",x"28",x"FC",x"B0",x"E9",
x"A2",x"25",x"20",x"82",x"F7",x"85",x"E0",x"20",
x"04",x"F8",x"60",x"A2",x"20",x"A9",x"16",x"20",
x"66",x"F7",x"CA",x"10",x"FA",x"A9",x"2A",x"20",
x"66",x"F7",x"60",x"A2",x"00",x"20",x"C7",x"FF",
x"C9",x"16",x"D0",x"03",x"E8",x"D0",x"F6",x"C9",
x"2A",x"D0",x"F0",x"E0",x"09",x"90",x"EC",x"60",
x"A2",x"00",x"BD",x"34",x"02",x"C9",x"2A",x"F0",
x"0C",x"DD",x"3A",x"02",x"F0",x"02",x"38",x"60",
x"E8",x"E0",x"06",x"90",x"ED",x"18",x"60",x"A2",
x"00",x"20",x"C7",x"FF",x"9D",x"3A",x"02",x"E8",
x"E0",x"06",x"90",x"F5",x"60",x"20",x"8B",x"FC",
x"AA",x"20",x"1B",x"FA",x"F0",x"1A",x"C9",x"2A",
x"D0",x"05",x"9D",x"34",x"02",x"D0",x"11",x"C9",
x"20",x"08",x"20",x"69",x"FF",x"28",x"90",x"E9",
x"9D",x"34",x"02",x"E8",x"E0",x"06",x"D0",x"E1",
x"86",x"E2",x"60",x"A2",x"2F",x"20",x"82",x"F7",
x"AA",x"BD",x"34",x"02",x"20",x"69",x"FF",x"20",
x"66",x"F7",x"E8",x"E0",x"06",x"90",x"F2",x"20",
x"04",x"F8",x"60",x"A2",x"0B",x"A9",x"00",x"9D",
x"34",x"02",x"CA",x"10",x"FA",x"60",x"20",x"8B",
x"FC",x"AA",x"B5",x"14",x"F0",x"0D",x"E8",x"B5",
x"14",x"F0",x"08",x"9D",x"33",x"02",x"E8",x"E0",
x"07",x"D0",x"F4",x"86",x"E2",x"A9",x"61",x"85",
x"13",x"60",x"20",x"32",x"F7",x"20",x"7B",x"FB",
x"20",x"03",x"FC",x"20",x"73",x"FC",x"60",x"20",
x"4D",x"FC",x"20",x"13",x"F8",x"20",x"D5",x"F9",
x"E0",x"02",x"F0",x"13",x"20",x"F0",x"F8",x"4C",
x"BF",x"FC",x"00",x"9D",x"34",x"C9",x"1C",x"F0",
x"03",x"4C",x"74",x"A3",x"4C",x"59",x"A3",x"20",
x"38",x"FD",x"20",x"B2",x"FC",x"A2",x"03",x"B5",
x"FC",x"20",x"66",x"F7",x"CA",x"10",x"F8",x"A0",
x"00",x"B1",x"FC",x"20",x"66",x"F7",x"20",x"33",
x"FF",x"90",x"F4",x"B0",x"35",x"20",x"4D",x"FC",
x"20",x"13",x"F8",x"20",x"D5",x"F9",x"C6",x"E0",
x"20",x"D6",x"FB",x"A2",x"03",x"20",x"C7",x"FF",
x"95",x"FC",x"CA",x"10",x"F8",x"A6",x"E1",x"F0",
x"0D",x"20",x"42",x"FD",x"A2",x"04",x"20",x"42",
x"FB",x"A2",x"01",x"20",x"3A",x"FD",x"A0",x"00",
x"20",x"C7",x"FF",x"91",x"FC",x"20",x"33",x"FF",
x"90",x"F4",x"20",x"3D",x"F7",x"4C",x"EA",x"F8",
x"A2",x"03",x"B5",x"FA",x"95",x"FC",x"CA",x"10",
x"F9",x"60",x"38",x"A5",x"FE",x"E5",x"FC",x"85",
x"F8",x"A5",x"FF",x"E5",x"FD",x"85",x"F9",x"60",
x"20",x"79",x"FD",x"A2",x"04",x"20",x"8B",x"FB",
x"A2",x"01",x"20",x"71",x"FD",x"A0",x"00",x"20",
x"C7",x"FF",x"91",x"FC",x"20",x"33",x"FF",x"90",
x"F4",x"20",x"84",x"F7",x"4C",x"31",x"F9",x"A2",
x"03",x"B5",x"FA",x"95",x"FC",x"CA",x"10",x"F9",
x"60",x"38",x"A5",x"FE",x"E5",x"FC",x"85",x"F8",
x"A5",x"FF",x"E5",x"FD",x"85",x"F9",x"60",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"A2",x"28",x"9A",x"D8",x"20",x"A2",x"F0",x"A9",
x"00",x"85",x"FC",x"85",x"FD",x"A8",x"F0",x"2E",
x"20",x"34",x"F8",x"29",x"7F",x"C9",x"2F",x"F0",
x"35",x"C9",x"47",x"F0",x"2E",x"C9",x"4C",x"F0",
x"65",x"C9",x"58",x"D0",x"0A",x"A9",x"FE",x"48",
x"A9",x"25",x"48",x"08",x"4C",x"49",x"F8",x"20",
x"CC",x"F7",x"30",x"DC",x"A2",x"02",x"20",x"25",
x"F8",x"A9",x"1A",x"20",x"D3",x"F0",x"B1",x"FC",
x"85",x"FA",x"20",x"E5",x"F7",x"20",x"04",x"F8",
x"4C",x"10",x"FE",x"6C",x"FC",x"00",x"20",x"34",
x"F8",x"29",x"7F",x"C9",x"2E",x"F0",x"B9",x"C9",
x"0D",x"D0",x"0F",x"E6",x"FC",x"D0",x"02",x"E6",
x"FD",x"A0",x"00",x"B1",x"FC",x"85",x"FA",x"4C",
x"7D",x"FE",x"20",x"CC",x"F7",x"30",x"DF",x"A2",
x"00",x"20",x"25",x"F8",x"A5",x"FA",x"91",x"FC",
x"A9",x"1A",x"20",x"D3",x"F0",x"20",x"E5",x"F7",
x"20",x"04",x"F8",x"4C",x"4E",x"FE",x"85",x"E0",
x"F0",x"C4",x"4C",x"C2",x"FF",x"50",x"3B",x"2F",
x"20",x"5A",x"41",x"51",x"2C",x"4D",x"4E",x"42",
x"56",x"43",x"58",x"4B",x"4A",x"48",x"47",x"46",
x"44",x"53",x"49",x"55",x"59",x"54",x"52",x"45",
x"57",x"00",x"00",x"0D",x"0A",x"4F",x"4C",x"2E",
x"00",x"0E",x"2D",x"3A",x"30",x"39",x"38",x"37",
x"36",x"35",x"34",x"33",x"32",x"31",x"54",x"B2",
x"13",x"75",x"80",x"C9",x"A3",x"B8",x"DB",x"06",
x"2D",x"C6",x"CC",x"97",x"BB",x"9A",x"16",x"1D",
x"03",x"0A",x"C2",x"0E",x"41",x"A0",x"79",x"D5",
x"00",x"45",x"00",x"00",x"32",x"88",x"3F",x"BF",
x"94",x"00",x"65",x"A9",x"AC",x"A6",x"B5",x"21",
x"61",x"6D",x"7D",x"26",x"38",x"4D",x"49",x"A9",
x"2A",x"8D",x"01",x"88",x"A9",x"FF",x"8D",x"00",
x"88",x"A9",x"2E",x"8D",x"01",x"88",x"A9",x"2C",
x"8D",x"03",x"88",x"60",x"48",x"AD",x"01",x"88",
x"09",x"04",x"8D",x"01",x"88",x"68",x"8D",x"00",
x"88",x"AD",x"02",x"88",x"4A",x"B0",x"0B",x"EA",
x"EA",x"EA",x"2C",x"02",x"88",x"30",x"FB",x"AD",
x"00",x"88",x"60",x"A2",x"00",x"BD",x"3A",x"02",
x"F0",x"08",x"20",x"69",x"FF",x"E8",x"E0",x"06",
x"D0",x"F3",x"60",x"E6",x"FC",x"D0",x"02",x"E6",
x"FD",x"A5",x"FC",x"C5",x"FE",x"D0",x"08",x"A5",
x"FD",x"C5",x"FF",x"D0",x"02",x"38",x"60",x"18",
x"60",x"09",x"08",x"01",x"0C",x"1A",x"1E",x"0A",
x"0E",x"8A",x"48",x"A2",x"0A",x"20",x"56",x"F7",
x"68",x"AA",x"68",x"60",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"20",x"EE",x"FF",x"48",x"2C",x"4E",x"02",
x"10",x"05",x"68",x"48",x"20",x"04",x"FF",x"2C",
x"05",x"02",x"10",x"09",x"68",x"48",x"20",x"5F",
x"F7",x"C9",x"0D",x"F0",x"CC",x"68",x"60",x"AA",
x"AA",x"AA",x"AA",x"4C",x"89",x"FB",x"AA",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"4C",x"50",
x"FB",x"AA",x"AD",x"12",x"02",x"D0",x"19",x"A9",
x"FE",x"8D",x"00",x"DF",x"2C",x"00",x"DF",x"70",
x"0F",x"A9",x"FB",x"8D",x"00",x"DF",x"2C",x"00",
x"DF",x"70",x"05",x"A9",x"03",x"4C",x"36",x"A6",
x"60",x"2C",x"2C",x"03",x"02",x"30",x"03",x"4C",
x"F0",x"F2",x"20",x"3E",x"F8",x"F0",x"0A",x"AD",
x"00",x"E0",x"4A",x"90",x"F5",x"AD",x"01",x"E0",
x"60",x"20",x"46",x"F7",x"4C",x"F0",x"F2",x"C2",
x"C0",x"A8",x"CE",x"10",x"DA",x"14",x"D8",x"AA",
x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",
x"AA",x"AA",x"AA",x"6C",x"18",x"02",x"6C",x"1A",
x"02",x"6C",x"1C",x"02",x"6C",x"1E",x"02",x"6C",
x"20",x"02",x"2E",x"02",x"00",x"F0",x"49",x"F8"
);
begin
process (address)
begin
	q <= romdata (to_integer(unsigned(address)));
end process;
end behavior;

